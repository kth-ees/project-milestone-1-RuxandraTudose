module alu #(
  BW = 16 // bitwidth
  ) (
  input  logic unsigned [BW-1:0] in_a,
  input  logic unsigned [BW-1:0] in_b,
  input  logic             [3:0] opcode,
  output logic unsigned [BW-1:0] out,
  output logic             [2:0] flags // {overflow, negative, zero}
  );

  //describe the ALU operations acording to the table
  always_comb begin
	out = '0; //output rule
	case(opcode) 
		3'd0: out = in_a + in_b;
		3'd1: out = in_a - in_b;
		3'd2: out = in_a && in_b;
		3'd3: out = in_a || in_b;
		3'd4: out = in_a ^ in_b;
		3'd5: out = in_a + 1;
		3'd6: out = in_a;
		3'd7: out = in_b;
		default: out = '0;
	endcase
  end

   //describe the behaviour of the flags
   always_comb begin
	flags = 3'b000; //output rule 
	
	//condition for addition overflow
	//the sum of two numbers with the same sign should not result in a number of opposite sign
	if(opcode == 3'b000 && ((in_a[BW-1] & in_b[BW-1] & ~out[BW-1]) |
				(~in_a[BW-1] & ~in_b[BW-1] & out[BW-1]))) begin
		flags[2] = 1'b1;
	end
	
	//condition for subtraction overflow
	//if A and out have different signs and A and B have different signs before subtraction => overflow
	//e.g : 3 - (-5) = 8 (1000 - which is interpreted as -8)
	else if(opcode == 3'b001 && ((in_a[BW-1] & ~in_b[BW-1] & ~out[BW-1]) |
				(~in_a[BW-1] & in_b[BW-1] & out[BW-1]))) begin
		 
		flags[2] = 1'b1;
	end else 
		flags[2] = 1'b0;
	
	flags[1] = out[BW-1]; //negative flag
	flags[0] = ~|out; //zero flag - apply nor on the bits of 'out' 

   end

endmodule

